
module decoder_4to16(

    input [3:0]a,
    input enable,
    output [15:0]d

    );

