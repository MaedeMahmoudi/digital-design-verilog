
module tb_ring_counter;
    