
module half( sum , ca)